module MasterController(
    
)
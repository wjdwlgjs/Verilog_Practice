module AlteraClock(
    // buttons and switches
    input key1_i,
    input key2_i,
    input key3_i,
    input set_switch_i,
)